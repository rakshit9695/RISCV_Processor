// Program Counter (32-bit) – increments +4 or branches
module PC(
    input  logic        clk,
    input  logic        rst,
    input  logic [31:0] pc_next,
    output logic [31:0] pc
);
    always_ff @(posedge clk or posedge rst) begin
        if (rst) pc <= 32'h0000_0000;
        else     pc <= pc_next;
    end
endmodule
